//------------------------------------------------------------------------------
//Verification Engineer: Rajkumar Raval
//Company Name: Personal Project.
//File Description: This file contains the WB agent package in which all the class based components of the 
//WB agent has been included  
//This class instantiates the agent and subscriber.
//License: Released under Creative Commons Attribution - BY
//------------------------------------------------------------------------------

package wb_agent_pkg;

`include "ovm_macros.svh"
import ovm_pkg::*;


`include "ovm_wb_transaction.svh"
`include "ovm_wb_sequence.svh"
`include "ovm_wb_sequencer.svh"
`include "ovm_wb_master_driver.svh"
`include "ovm_wb_monitor.svh"
`include "ovm_wb_agent.svh"
`include "ovm_wb_subscriber.svh"

endpackage
